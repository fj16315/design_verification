-- *****************************************************************
-- Specman Elite VHDL stubs file: /home/fj16315/linux/Documents/3rd_Year/Design_Verification/Assignment_2/INCA_libs/irun.lnx8664.14.10.nc/specman.14.10.004-s/scratch/specman.vhd
-- Topmost e module: calc1_sn_env.e
-- Generated using seed = 1
-- Generated using separator : ':' 
-- Date: Mon Dec 10 13:29:43 2018
-- Specman Elite version: 14.10.004-s
-- *****************************************************************

entity SPECMAN_FMI is
     generic (
ncrun : string := "ncrun"
     );
end SPECMAN_FMI;
architecture fmi_stub of SPECMAN_FMI is
 attribute FOREIGN of fmi_stub: architecture is "SN_C_MODEL:SN_SPECMAN";
begin
end fmi_stub;


entity SPECMAN_VHPI is
end SPECMAN_VHPI;
architecture vhpi_stub of SPECMAN_VHPI is
 attribute FOREIGN of vhpi_stub: architecture is "VHPIDIRECT libncvhdl_sn_boot: sn_vhpi_arch_elab sn_vhpi_arch_exec";
begin
end vhpi_stub;


library IEEE;
use IEEE.std_logic_1164.all;

entity  specman_wave_vhdl is
end specman_wave_vhdl;
architecture arch of specman_wave_vhdl is 
  constant sn_integer_num: integer := 100;
  constant sn_boolean_num: integer := 100;
  constant sn_error_num:integer := 1;
  constant sn_error_len: integer := 80;
  constant sn_message_num: integer := 3;
  constant sn_message_len: integer := 80;
  constant sn_string_num: integer := 200;
  constant sn_string_len: integer := 80;
  constant sn_event_num: integer := 0;
  type sn_intg_array is array (NATURAL range <>) of integer;
  subtype sn_error_string is string (1 to 80);
  subtype sn_msg_string is string (1 to 80);
  subtype sn_string is string (1 to 80);
  signal sn_intg1: integer;
  signal sn_intg2: integer;
  signal sn_intg3: integer;
  signal sn_intg4: integer;
  signal sn_intg5: integer;
  signal sn_intg6: integer;
  signal sn_intg7: integer;
  signal sn_intg8: integer;
  signal sn_intg9: integer;
  signal sn_intg10: integer;
  signal sn_intg11: integer;
  signal sn_intg12: integer;
  signal sn_intg13: integer;
  signal sn_intg14: integer;
  signal sn_intg15: integer;
  signal sn_intg16: integer;
  signal sn_intg17: integer;
  signal sn_intg18: integer;
  signal sn_intg19: integer;
  signal sn_intg20: integer;
  signal sn_intg21: integer;
  signal sn_intg22: integer;
  signal sn_intg23: integer;
  signal sn_intg24: integer;
  signal sn_intg25: integer;
  signal sn_intg26: integer;
  signal sn_intg27: integer;
  signal sn_intg28: integer;
  signal sn_intg29: integer;
  signal sn_intg30: integer;
  signal sn_intg31: integer;
  signal sn_intg32: integer;
  signal sn_intg33: integer;
  signal sn_intg34: integer;
  signal sn_intg35: integer;
  signal sn_intg36: integer;
  signal sn_intg37: integer;
  signal sn_intg38: integer;
  signal sn_intg39: integer;
  signal sn_intg40: integer;
  signal sn_intg41: integer;
  signal sn_intg42: integer;
  signal sn_intg43: integer;
  signal sn_intg44: integer;
  signal sn_intg45: integer;
  signal sn_intg46: integer;
  signal sn_intg47: integer;
  signal sn_intg48: integer;
  signal sn_intg49: integer;
  signal sn_intg50: integer;
  signal sn_intg51: integer;
  signal sn_intg52: integer;
  signal sn_intg53: integer;
  signal sn_intg54: integer;
  signal sn_intg55: integer;
  signal sn_intg56: integer;
  signal sn_intg57: integer;
  signal sn_intg58: integer;
  signal sn_intg59: integer;
  signal sn_intg60: integer;
  signal sn_intg61: integer;
  signal sn_intg62: integer;
  signal sn_intg63: integer;
  signal sn_intg64: integer;
  signal sn_intg65: integer;
  signal sn_intg66: integer;
  signal sn_intg67: integer;
  signal sn_intg68: integer;
  signal sn_intg69: integer;
  signal sn_intg70: integer;
  signal sn_intg71: integer;
  signal sn_intg72: integer;
  signal sn_intg73: integer;
  signal sn_intg74: integer;
  signal sn_intg75: integer;
  signal sn_intg76: integer;
  signal sn_intg77: integer;
  signal sn_intg78: integer;
  signal sn_intg79: integer;
  signal sn_intg80: integer;
  signal sn_intg81: integer;
  signal sn_intg82: integer;
  signal sn_intg83: integer;
  signal sn_intg84: integer;
  signal sn_intg85: integer;
  signal sn_intg86: integer;
  signal sn_intg87: integer;
  signal sn_intg88: integer;
  signal sn_intg89: integer;
  signal sn_intg90: integer;
  signal sn_intg91: integer;
  signal sn_intg92: integer;
  signal sn_intg93: integer;
  signal sn_intg94: integer;
  signal sn_intg95: integer;
  signal sn_intg96: integer;
  signal sn_intg97: integer;
  signal sn_intg98: integer;
  signal sn_intg99: integer;
  signal sn_intg100: integer;
  signal sn_bool1: std_ulogic;
  signal sn_bool2: std_ulogic;
  signal sn_bool3: std_ulogic;
  signal sn_bool4: std_ulogic;
  signal sn_bool5: std_ulogic;
  signal sn_bool6: std_ulogic;
  signal sn_bool7: std_ulogic;
  signal sn_bool8: std_ulogic;
  signal sn_bool9: std_ulogic;
  signal sn_bool10: std_ulogic;
  signal sn_bool11: std_ulogic;
  signal sn_bool12: std_ulogic;
  signal sn_bool13: std_ulogic;
  signal sn_bool14: std_ulogic;
  signal sn_bool15: std_ulogic;
  signal sn_bool16: std_ulogic;
  signal sn_bool17: std_ulogic;
  signal sn_bool18: std_ulogic;
  signal sn_bool19: std_ulogic;
  signal sn_bool20: std_ulogic;
  signal sn_bool21: std_ulogic;
  signal sn_bool22: std_ulogic;
  signal sn_bool23: std_ulogic;
  signal sn_bool24: std_ulogic;
  signal sn_bool25: std_ulogic;
  signal sn_bool26: std_ulogic;
  signal sn_bool27: std_ulogic;
  signal sn_bool28: std_ulogic;
  signal sn_bool29: std_ulogic;
  signal sn_bool30: std_ulogic;
  signal sn_bool31: std_ulogic;
  signal sn_bool32: std_ulogic;
  signal sn_bool33: std_ulogic;
  signal sn_bool34: std_ulogic;
  signal sn_bool35: std_ulogic;
  signal sn_bool36: std_ulogic;
  signal sn_bool37: std_ulogic;
  signal sn_bool38: std_ulogic;
  signal sn_bool39: std_ulogic;
  signal sn_bool40: std_ulogic;
  signal sn_bool41: std_ulogic;
  signal sn_bool42: std_ulogic;
  signal sn_bool43: std_ulogic;
  signal sn_bool44: std_ulogic;
  signal sn_bool45: std_ulogic;
  signal sn_bool46: std_ulogic;
  signal sn_bool47: std_ulogic;
  signal sn_bool48: std_ulogic;
  signal sn_bool49: std_ulogic;
  signal sn_bool50: std_ulogic;
  signal sn_bool51: std_ulogic;
  signal sn_bool52: std_ulogic;
  signal sn_bool53: std_ulogic;
  signal sn_bool54: std_ulogic;
  signal sn_bool55: std_ulogic;
  signal sn_bool56: std_ulogic;
  signal sn_bool57: std_ulogic;
  signal sn_bool58: std_ulogic;
  signal sn_bool59: std_ulogic;
  signal sn_bool60: std_ulogic;
  signal sn_bool61: std_ulogic;
  signal sn_bool62: std_ulogic;
  signal sn_bool63: std_ulogic;
  signal sn_bool64: std_ulogic;
  signal sn_bool65: std_ulogic;
  signal sn_bool66: std_ulogic;
  signal sn_bool67: std_ulogic;
  signal sn_bool68: std_ulogic;
  signal sn_bool69: std_ulogic;
  signal sn_bool70: std_ulogic;
  signal sn_bool71: std_ulogic;
  signal sn_bool72: std_ulogic;
  signal sn_bool73: std_ulogic;
  signal sn_bool74: std_ulogic;
  signal sn_bool75: std_ulogic;
  signal sn_bool76: std_ulogic;
  signal sn_bool77: std_ulogic;
  signal sn_bool78: std_ulogic;
  signal sn_bool79: std_ulogic;
  signal sn_bool80: std_ulogic;
  signal sn_bool81: std_ulogic;
  signal sn_bool82: std_ulogic;
  signal sn_bool83: std_ulogic;
  signal sn_bool84: std_ulogic;
  signal sn_bool85: std_ulogic;
  signal sn_bool86: std_ulogic;
  signal sn_bool87: std_ulogic;
  signal sn_bool88: std_ulogic;
  signal sn_bool89: std_ulogic;
  signal sn_bool90: std_ulogic;
  signal sn_bool91: std_ulogic;
  signal sn_bool92: std_ulogic;
  signal sn_bool93: std_ulogic;
  signal sn_bool94: std_ulogic;
  signal sn_bool95: std_ulogic;
  signal sn_bool96: std_ulogic;
  signal sn_bool97: std_ulogic;
  signal sn_bool98: std_ulogic;
  signal sn_bool99: std_ulogic;
  signal sn_bool100: std_ulogic;
  signal sn_err_str1: sn_error_string := (others => ' ');
  signal sn_msg_str1: sn_msg_string := (others => ' ');
  signal sn_msg_str2: sn_msg_string := (others => ' ');
  signal sn_msg_str3: sn_msg_string := (others => ' ');
  signal sn_str1: sn_string := (others => ' ');
  signal sn_str2: sn_string := (others => ' ');
  signal sn_str3: sn_string := (others => ' ');
  signal sn_str4: sn_string := (others => ' ');
  signal sn_str5: sn_string := (others => ' ');
  signal sn_str6: sn_string := (others => ' ');
  signal sn_str7: sn_string := (others => ' ');
  signal sn_str8: sn_string := (others => ' ');
  signal sn_str9: sn_string := (others => ' ');
  signal sn_str10: sn_string := (others => ' ');
  signal sn_str11: sn_string := (others => ' ');
  signal sn_str12: sn_string := (others => ' ');
  signal sn_str13: sn_string := (others => ' ');
  signal sn_str14: sn_string := (others => ' ');
  signal sn_str15: sn_string := (others => ' ');
  signal sn_str16: sn_string := (others => ' ');
  signal sn_str17: sn_string := (others => ' ');
  signal sn_str18: sn_string := (others => ' ');
  signal sn_str19: sn_string := (others => ' ');
  signal sn_str20: sn_string := (others => ' ');
  signal sn_str21: sn_string := (others => ' ');
  signal sn_str22: sn_string := (others => ' ');
  signal sn_str23: sn_string := (others => ' ');
  signal sn_str24: sn_string := (others => ' ');
  signal sn_str25: sn_string := (others => ' ');
  signal sn_str26: sn_string := (others => ' ');
  signal sn_str27: sn_string := (others => ' ');
  signal sn_str28: sn_string := (others => ' ');
  signal sn_str29: sn_string := (others => ' ');
  signal sn_str30: sn_string := (others => ' ');
  signal sn_str31: sn_string := (others => ' ');
  signal sn_str32: sn_string := (others => ' ');
  signal sn_str33: sn_string := (others => ' ');
  signal sn_str34: sn_string := (others => ' ');
  signal sn_str35: sn_string := (others => ' ');
  signal sn_str36: sn_string := (others => ' ');
  signal sn_str37: sn_string := (others => ' ');
  signal sn_str38: sn_string := (others => ' ');
  signal sn_str39: sn_string := (others => ' ');
  signal sn_str40: sn_string := (others => ' ');
  signal sn_str41: sn_string := (others => ' ');
  signal sn_str42: sn_string := (others => ' ');
  signal sn_str43: sn_string := (others => ' ');
  signal sn_str44: sn_string := (others => ' ');
  signal sn_str45: sn_string := (others => ' ');
  signal sn_str46: sn_string := (others => ' ');
  signal sn_str47: sn_string := (others => ' ');
  signal sn_str48: sn_string := (others => ' ');
  signal sn_str49: sn_string := (others => ' ');
  signal sn_str50: sn_string := (others => ' ');
  signal sn_str51: sn_string := (others => ' ');
  signal sn_str52: sn_string := (others => ' ');
  signal sn_str53: sn_string := (others => ' ');
  signal sn_str54: sn_string := (others => ' ');
  signal sn_str55: sn_string := (others => ' ');
  signal sn_str56: sn_string := (others => ' ');
  signal sn_str57: sn_string := (others => ' ');
  signal sn_str58: sn_string := (others => ' ');
  signal sn_str59: sn_string := (others => ' ');
  signal sn_str60: sn_string := (others => ' ');
  signal sn_str61: sn_string := (others => ' ');
  signal sn_str62: sn_string := (others => ' ');
  signal sn_str63: sn_string := (others => ' ');
  signal sn_str64: sn_string := (others => ' ');
  signal sn_str65: sn_string := (others => ' ');
  signal sn_str66: sn_string := (others => ' ');
  signal sn_str67: sn_string := (others => ' ');
  signal sn_str68: sn_string := (others => ' ');
  signal sn_str69: sn_string := (others => ' ');
  signal sn_str70: sn_string := (others => ' ');
  signal sn_str71: sn_string := (others => ' ');
  signal sn_str72: sn_string := (others => ' ');
  signal sn_str73: sn_string := (others => ' ');
  signal sn_str74: sn_string := (others => ' ');
  signal sn_str75: sn_string := (others => ' ');
  signal sn_str76: sn_string := (others => ' ');
  signal sn_str77: sn_string := (others => ' ');
  signal sn_str78: sn_string := (others => ' ');
  signal sn_str79: sn_string := (others => ' ');
  signal sn_str80: sn_string := (others => ' ');
  signal sn_str81: sn_string := (others => ' ');
  signal sn_str82: sn_string := (others => ' ');
  signal sn_str83: sn_string := (others => ' ');
  signal sn_str84: sn_string := (others => ' ');
  signal sn_str85: sn_string := (others => ' ');
  signal sn_str86: sn_string := (others => ' ');
  signal sn_str87: sn_string := (others => ' ');
  signal sn_str88: sn_string := (others => ' ');
  signal sn_str89: sn_string := (others => ' ');
  signal sn_str90: sn_string := (others => ' ');
  signal sn_str91: sn_string := (others => ' ');
  signal sn_str92: sn_string := (others => ' ');
  signal sn_str93: sn_string := (others => ' ');
  signal sn_str94: sn_string := (others => ' ');
  signal sn_str95: sn_string := (others => ' ');
  signal sn_str96: sn_string := (others => ' ');
  signal sn_str97: sn_string := (others => ' ');
  signal sn_str98: sn_string := (others => ' ');
  signal sn_str99: sn_string := (others => ' ');
  signal sn_str100: sn_string := (others => ' ');
  signal sn_str101: sn_string := (others => ' ');
  signal sn_str102: sn_string := (others => ' ');
  signal sn_str103: sn_string := (others => ' ');
  signal sn_str104: sn_string := (others => ' ');
  signal sn_str105: sn_string := (others => ' ');
  signal sn_str106: sn_string := (others => ' ');
  signal sn_str107: sn_string := (others => ' ');
  signal sn_str108: sn_string := (others => ' ');
  signal sn_str109: sn_string := (others => ' ');
  signal sn_str110: sn_string := (others => ' ');
  signal sn_str111: sn_string := (others => ' ');
  signal sn_str112: sn_string := (others => ' ');
  signal sn_str113: sn_string := (others => ' ');
  signal sn_str114: sn_string := (others => ' ');
  signal sn_str115: sn_string := (others => ' ');
  signal sn_str116: sn_string := (others => ' ');
  signal sn_str117: sn_string := (others => ' ');
  signal sn_str118: sn_string := (others => ' ');
  signal sn_str119: sn_string := (others => ' ');
  signal sn_str120: sn_string := (others => ' ');
  signal sn_str121: sn_string := (others => ' ');
  signal sn_str122: sn_string := (others => ' ');
  signal sn_str123: sn_string := (others => ' ');
  signal sn_str124: sn_string := (others => ' ');
  signal sn_str125: sn_string := (others => ' ');
  signal sn_str126: sn_string := (others => ' ');
  signal sn_str127: sn_string := (others => ' ');
  signal sn_str128: sn_string := (others => ' ');
  signal sn_str129: sn_string := (others => ' ');
  signal sn_str130: sn_string := (others => ' ');
  signal sn_str131: sn_string := (others => ' ');
  signal sn_str132: sn_string := (others => ' ');
  signal sn_str133: sn_string := (others => ' ');
  signal sn_str134: sn_string := (others => ' ');
  signal sn_str135: sn_string := (others => ' ');
  signal sn_str136: sn_string := (others => ' ');
  signal sn_str137: sn_string := (others => ' ');
  signal sn_str138: sn_string := (others => ' ');
  signal sn_str139: sn_string := (others => ' ');
  signal sn_str140: sn_string := (others => ' ');
  signal sn_str141: sn_string := (others => ' ');
  signal sn_str142: sn_string := (others => ' ');
  signal sn_str143: sn_string := (others => ' ');
  signal sn_str144: sn_string := (others => ' ');
  signal sn_str145: sn_string := (others => ' ');
  signal sn_str146: sn_string := (others => ' ');
  signal sn_str147: sn_string := (others => ' ');
  signal sn_str148: sn_string := (others => ' ');
  signal sn_str149: sn_string := (others => ' ');
  signal sn_str150: sn_string := (others => ' ');
  signal sn_str151: sn_string := (others => ' ');
  signal sn_str152: sn_string := (others => ' ');
  signal sn_str153: sn_string := (others => ' ');
  signal sn_str154: sn_string := (others => ' ');
  signal sn_str155: sn_string := (others => ' ');
  signal sn_str156: sn_string := (others => ' ');
  signal sn_str157: sn_string := (others => ' ');
  signal sn_str158: sn_string := (others => ' ');
  signal sn_str159: sn_string := (others => ' ');
  signal sn_str160: sn_string := (others => ' ');
  signal sn_str161: sn_string := (others => ' ');
  signal sn_str162: sn_string := (others => ' ');
  signal sn_str163: sn_string := (others => ' ');
  signal sn_str164: sn_string := (others => ' ');
  signal sn_str165: sn_string := (others => ' ');
  signal sn_str166: sn_string := (others => ' ');
  signal sn_str167: sn_string := (others => ' ');
  signal sn_str168: sn_string := (others => ' ');
  signal sn_str169: sn_string := (others => ' ');
  signal sn_str170: sn_string := (others => ' ');
  signal sn_str171: sn_string := (others => ' ');
  signal sn_str172: sn_string := (others => ' ');
  signal sn_str173: sn_string := (others => ' ');
  signal sn_str174: sn_string := (others => ' ');
  signal sn_str175: sn_string := (others => ' ');
  signal sn_str176: sn_string := (others => ' ');
  signal sn_str177: sn_string := (others => ' ');
  signal sn_str178: sn_string := (others => ' ');
  signal sn_str179: sn_string := (others => ' ');
  signal sn_str180: sn_string := (others => ' ');
  signal sn_str181: sn_string := (others => ' ');
  signal sn_str182: sn_string := (others => ' ');
  signal sn_str183: sn_string := (others => ' ');
  signal sn_str184: sn_string := (others => ' ');
  signal sn_str185: sn_string := (others => ' ');
  signal sn_str186: sn_string := (others => ' ');
  signal sn_str187: sn_string := (others => ' ');
  signal sn_str188: sn_string := (others => ' ');
  signal sn_str189: sn_string := (others => ' ');
  signal sn_str190: sn_string := (others => ' ');
  signal sn_str191: sn_string := (others => ' ');
  signal sn_str192: sn_string := (others => ' ');
  signal sn_str193: sn_string := (others => ' ');
  signal sn_str194: sn_string := (others => ' ');
  signal sn_str195: sn_string := (others => ' ');
  signal sn_str196: sn_string := (others => ' ');
  signal sn_str197: sn_string := (others => ' ');
  signal sn_str198: sn_string := (others => ' ');
  signal sn_str199: sn_string := (others => ' ');
  signal sn_str200: sn_string := (others => ' ');
begin 
end arch;
  
  
   library IEEE; 

   use IEEE.std_logic_1164.all;

entity SPECMAN_REFERENCE is
end SPECMAN_REFERENCE;

architecture arch of SPECMAN_REFERENCE is

   component SN
   end component;

   for all: SN use entity work.SPECMAN_FMI(fmi_stub);

   component SN2
   end component;

   for all: SN2 use entity work.SPECMAN_VHPI(vhpi_stub);

   component SN_WAVE
   end component;

   for all: SN_WAVE use entity work.specman_wave_vhdl;

   --Specman stub attributes
   constant sn_version_id: integer := 0;
   constant sn_version_date: integer := 1310706;
   constant sn_use_wave: integer := 1;
   constant sn_port_unification : integer := 2; -- 1 for enabled, 2 for disabled
   constant sn_stub_elab: integer := 0;
   signal sn_control: integer := 0;
   signal sn_control_cb: integer := 0;
 begin
   sn_control_cb <= sn_control;
   SN_INST : SN;
   SN_INST2 : SN2;
   SN_WAVE_INST : SN_WAVE;
 end arch;

